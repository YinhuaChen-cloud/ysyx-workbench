module IDU(
  input  [31:0] io_inst,
  input         io_idu_to_exu_br_eq,
  input         io_idu_to_exu_br_lt,
  input         io_idu_to_exu_br_ltu,
  output [3:0]  io_idu_to_exu_pc_sel,
  output [1:0]  io_idu_to_exu_op1_sel,
  output [2:0]  io_idu_to_exu_op2_sel,
  output [3:0]  io_idu_to_exu_alu_op,
  output [1:0]  io_idu_to_exu_wb_sel,
  output        io_idu_to_exu_reg_wen,
  output [2:0]  io_idu_to_exu_mem_msk_type,
  output        io_idu_to_exu_alu_msk_type,
  output        io_isEbreak,
  output        io_inv_inst,
  output        io_isWriteMem
);
  wire [31:0] _decoded_signals_T = io_inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_1 = 32'h33 == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_3 = 32'h3b == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_5 = 32'h40000033 == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_7 = 32'h4000003b == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_9 = 32'h2000033 == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_11 = 32'h200003b == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_13 = 32'h200403b == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_15 = 32'h2005033 == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_17 = 32'h200503b == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_19 = 32'h200603b == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_21 = 32'h1033 == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_23 = 32'h103b == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_25 = 32'h503b == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_27 = 32'h4000503b == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_29 = 32'h7033 == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_31 = 32'h6033 == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_33 = 32'h4033 == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_35 = 32'h2033 == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_37 = 32'h3033 == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire [31:0] _decoded_signals_T_38 = io_inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_39 = 32'h3003 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_41 = 32'h2003 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_43 = 32'h6003 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_45 = 32'h1003 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_47 = 32'h5003 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_49 = 32'h3 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_51 = 32'h4003 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_53 = 32'h13 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_55 = 32'h1b == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire [31:0] _decoded_signals_T_56 = io_inst & 32'hfc00707f; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_57 = 32'h1013 == _decoded_signals_T_56; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_59 = 32'h101b == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_61 = 32'h5013 == _decoded_signals_T_56; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_63 = 32'h501b == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_65 = 32'h40005013 == _decoded_signals_T_56; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_67 = 32'h4000501b == _decoded_signals_T; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_69 = 32'h7013 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_71 = 32'h6013 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_73 = 32'h4013 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_75 = 32'h67 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_77 = 32'h3013 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_79 = 32'h3023 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_81 = 32'h2023 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_83 = 32'h1023 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_85 = 32'h23 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_87 = 32'h63 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_89 = 32'h1063 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_91 = 32'h5063 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_93 = 32'h7063 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_95 = 32'h4063 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_97 = 32'h6063 == _decoded_signals_T_38; // @[Lookup.scala 31:38]
  wire [31:0] _decoded_signals_T_98 = io_inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_99 = 32'h37 == _decoded_signals_T_98; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_101 = 32'h17 == _decoded_signals_T_98; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_103 = 32'h6f == _decoded_signals_T_98; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_105 = 32'h100073 == io_inst; // @[Lookup.scala 31:38]
  wire  _decoded_signals_T_136 = _decoded_signals_T_45 | (_decoded_signals_T_47 | (_decoded_signals_T_49 | (
    _decoded_signals_T_51 | (_decoded_signals_T_53 | (_decoded_signals_T_55 | (_decoded_signals_T_57 | (
    _decoded_signals_T_59 | (_decoded_signals_T_61 | (_decoded_signals_T_63 | (_decoded_signals_T_65 | (
    _decoded_signals_T_67 | (_decoded_signals_T_69 | (_decoded_signals_T_71 | (_decoded_signals_T_73 | (
    _decoded_signals_T_75 | (_decoded_signals_T_77 | (_decoded_signals_T_79 | (_decoded_signals_T_81 | (
    _decoded_signals_T_83 | (_decoded_signals_T_85 | (_decoded_signals_T_87 | (_decoded_signals_T_89 | (
    _decoded_signals_T_91 | (_decoded_signals_T_93 | (_decoded_signals_T_95 | (_decoded_signals_T_97 | (
    _decoded_signals_T_99 | (_decoded_signals_T_101 | (_decoded_signals_T_103 | _decoded_signals_T_105))))))))))))))))))
    ))))))))))); // @[Lookup.scala 34:39]
  wire  decoded_signals_0 = _decoded_signals_T_1 | (_decoded_signals_T_3 | (_decoded_signals_T_5 | (_decoded_signals_T_7
     | (_decoded_signals_T_9 | (_decoded_signals_T_11 | (_decoded_signals_T_13 | (_decoded_signals_T_15 | (
    _decoded_signals_T_17 | (_decoded_signals_T_19 | (_decoded_signals_T_21 | (_decoded_signals_T_23 | (
    _decoded_signals_T_25 | (_decoded_signals_T_27 | (_decoded_signals_T_29 | (_decoded_signals_T_31 | (
    _decoded_signals_T_33 | (_decoded_signals_T_35 | (_decoded_signals_T_37 | (_decoded_signals_T_39 | (
    _decoded_signals_T_41 | (_decoded_signals_T_43 | _decoded_signals_T_136))))))))))))))))))))); // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_159 = _decoded_signals_T_103 ? 4'h7 : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_160 = _decoded_signals_T_101 ? 4'h0 : _decoded_signals_T_159; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_161 = _decoded_signals_T_99 ? 4'h0 : _decoded_signals_T_160; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_162 = _decoded_signals_T_97 ? 4'h6 : _decoded_signals_T_161; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_163 = _decoded_signals_T_95 ? 4'h5 : _decoded_signals_T_162; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_164 = _decoded_signals_T_93 ? 4'h4 : _decoded_signals_T_163; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_165 = _decoded_signals_T_91 ? 4'h3 : _decoded_signals_T_164; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_166 = _decoded_signals_T_89 ? 4'h1 : _decoded_signals_T_165; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_167 = _decoded_signals_T_87 ? 4'h2 : _decoded_signals_T_166; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_168 = _decoded_signals_T_85 ? 4'h0 : _decoded_signals_T_167; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_169 = _decoded_signals_T_83 ? 4'h0 : _decoded_signals_T_168; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_170 = _decoded_signals_T_81 ? 4'h0 : _decoded_signals_T_169; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_171 = _decoded_signals_T_79 ? 4'h0 : _decoded_signals_T_170; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_172 = _decoded_signals_T_77 ? 4'h0 : _decoded_signals_T_171; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_173 = _decoded_signals_T_75 ? 4'h8 : _decoded_signals_T_172; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_174 = _decoded_signals_T_73 ? 4'h0 : _decoded_signals_T_173; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_175 = _decoded_signals_T_71 ? 4'h0 : _decoded_signals_T_174; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_176 = _decoded_signals_T_69 ? 4'h0 : _decoded_signals_T_175; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_177 = _decoded_signals_T_67 ? 4'h0 : _decoded_signals_T_176; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_178 = _decoded_signals_T_65 ? 4'h0 : _decoded_signals_T_177; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_179 = _decoded_signals_T_63 ? 4'h0 : _decoded_signals_T_178; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_180 = _decoded_signals_T_61 ? 4'h0 : _decoded_signals_T_179; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_181 = _decoded_signals_T_59 ? 4'h0 : _decoded_signals_T_180; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_182 = _decoded_signals_T_57 ? 4'h0 : _decoded_signals_T_181; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_183 = _decoded_signals_T_55 ? 4'h0 : _decoded_signals_T_182; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_184 = _decoded_signals_T_53 ? 4'h0 : _decoded_signals_T_183; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_185 = _decoded_signals_T_51 ? 4'h0 : _decoded_signals_T_184; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_186 = _decoded_signals_T_49 ? 4'h0 : _decoded_signals_T_185; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_187 = _decoded_signals_T_47 ? 4'h0 : _decoded_signals_T_186; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_188 = _decoded_signals_T_45 ? 4'h0 : _decoded_signals_T_187; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_189 = _decoded_signals_T_43 ? 4'h0 : _decoded_signals_T_188; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_190 = _decoded_signals_T_41 ? 4'h0 : _decoded_signals_T_189; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_191 = _decoded_signals_T_39 ? 4'h0 : _decoded_signals_T_190; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_192 = _decoded_signals_T_37 ? 4'h0 : _decoded_signals_T_191; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_193 = _decoded_signals_T_35 ? 4'h0 : _decoded_signals_T_192; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_194 = _decoded_signals_T_33 ? 4'h0 : _decoded_signals_T_193; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_195 = _decoded_signals_T_31 ? 4'h0 : _decoded_signals_T_194; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_196 = _decoded_signals_T_29 ? 4'h0 : _decoded_signals_T_195; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_197 = _decoded_signals_T_27 ? 4'h0 : _decoded_signals_T_196; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_198 = _decoded_signals_T_25 ? 4'h0 : _decoded_signals_T_197; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_199 = _decoded_signals_T_23 ? 4'h0 : _decoded_signals_T_198; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_200 = _decoded_signals_T_21 ? 4'h0 : _decoded_signals_T_199; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_201 = _decoded_signals_T_19 ? 4'h0 : _decoded_signals_T_200; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_202 = _decoded_signals_T_17 ? 4'h0 : _decoded_signals_T_201; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_203 = _decoded_signals_T_15 ? 4'h0 : _decoded_signals_T_202; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_204 = _decoded_signals_T_13 ? 4'h0 : _decoded_signals_T_203; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_205 = _decoded_signals_T_11 ? 4'h0 : _decoded_signals_T_204; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_206 = _decoded_signals_T_9 ? 4'h0 : _decoded_signals_T_205; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_207 = _decoded_signals_T_7 ? 4'h0 : _decoded_signals_T_206; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_208 = _decoded_signals_T_5 ? 4'h0 : _decoded_signals_T_207; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_209 = _decoded_signals_T_3 ? 4'h0 : _decoded_signals_T_208; // @[Lookup.scala 34:39]
  wire [3:0] br_type = _decoded_signals_T_1 ? 4'h0 : _decoded_signals_T_209; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_212 = _decoded_signals_T_101 ? 2'h2 : 2'h0; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_213 = _decoded_signals_T_99 ? 2'h2 : _decoded_signals_T_212; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_214 = _decoded_signals_T_97 ? 2'h0 : _decoded_signals_T_213; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_215 = _decoded_signals_T_95 ? 2'h0 : _decoded_signals_T_214; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_216 = _decoded_signals_T_93 ? 2'h0 : _decoded_signals_T_215; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_217 = _decoded_signals_T_91 ? 2'h0 : _decoded_signals_T_216; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_218 = _decoded_signals_T_89 ? 2'h0 : _decoded_signals_T_217; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_219 = _decoded_signals_T_87 ? 2'h0 : _decoded_signals_T_218; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_220 = _decoded_signals_T_85 ? 2'h1 : _decoded_signals_T_219; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_221 = _decoded_signals_T_83 ? 2'h1 : _decoded_signals_T_220; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_222 = _decoded_signals_T_81 ? 2'h1 : _decoded_signals_T_221; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_223 = _decoded_signals_T_79 ? 2'h1 : _decoded_signals_T_222; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_224 = _decoded_signals_T_77 ? 2'h1 : _decoded_signals_T_223; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_225 = _decoded_signals_T_75 ? 2'h1 : _decoded_signals_T_224; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_226 = _decoded_signals_T_73 ? 2'h1 : _decoded_signals_T_225; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_227 = _decoded_signals_T_71 ? 2'h1 : _decoded_signals_T_226; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_228 = _decoded_signals_T_69 ? 2'h1 : _decoded_signals_T_227; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_229 = _decoded_signals_T_67 ? 2'h1 : _decoded_signals_T_228; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_230 = _decoded_signals_T_65 ? 2'h1 : _decoded_signals_T_229; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_231 = _decoded_signals_T_63 ? 2'h1 : _decoded_signals_T_230; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_232 = _decoded_signals_T_61 ? 2'h1 : _decoded_signals_T_231; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_233 = _decoded_signals_T_59 ? 2'h1 : _decoded_signals_T_232; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_234 = _decoded_signals_T_57 ? 2'h1 : _decoded_signals_T_233; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_235 = _decoded_signals_T_55 ? 2'h1 : _decoded_signals_T_234; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_236 = _decoded_signals_T_53 ? 2'h1 : _decoded_signals_T_235; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_237 = _decoded_signals_T_51 ? 2'h1 : _decoded_signals_T_236; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_238 = _decoded_signals_T_49 ? 2'h1 : _decoded_signals_T_237; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_239 = _decoded_signals_T_47 ? 2'h1 : _decoded_signals_T_238; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_240 = _decoded_signals_T_45 ? 2'h1 : _decoded_signals_T_239; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_241 = _decoded_signals_T_43 ? 2'h1 : _decoded_signals_T_240; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_242 = _decoded_signals_T_41 ? 2'h1 : _decoded_signals_T_241; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_243 = _decoded_signals_T_39 ? 2'h1 : _decoded_signals_T_242; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_244 = _decoded_signals_T_37 ? 2'h1 : _decoded_signals_T_243; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_245 = _decoded_signals_T_35 ? 2'h1 : _decoded_signals_T_244; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_246 = _decoded_signals_T_33 ? 2'h1 : _decoded_signals_T_245; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_247 = _decoded_signals_T_31 ? 2'h1 : _decoded_signals_T_246; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_248 = _decoded_signals_T_29 ? 2'h1 : _decoded_signals_T_247; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_249 = _decoded_signals_T_27 ? 2'h1 : _decoded_signals_T_248; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_250 = _decoded_signals_T_25 ? 2'h1 : _decoded_signals_T_249; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_251 = _decoded_signals_T_23 ? 2'h1 : _decoded_signals_T_250; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_252 = _decoded_signals_T_21 ? 2'h1 : _decoded_signals_T_251; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_253 = _decoded_signals_T_19 ? 2'h1 : _decoded_signals_T_252; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_254 = _decoded_signals_T_17 ? 2'h1 : _decoded_signals_T_253; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_255 = _decoded_signals_T_15 ? 2'h1 : _decoded_signals_T_254; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_256 = _decoded_signals_T_13 ? 2'h1 : _decoded_signals_T_255; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_257 = _decoded_signals_T_11 ? 2'h1 : _decoded_signals_T_256; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_258 = _decoded_signals_T_9 ? 2'h1 : _decoded_signals_T_257; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_259 = _decoded_signals_T_7 ? 2'h1 : _decoded_signals_T_258; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_260 = _decoded_signals_T_5 ? 2'h1 : _decoded_signals_T_259; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_261 = _decoded_signals_T_3 ? 2'h1 : _decoded_signals_T_260; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_264 = _decoded_signals_T_101 ? 3'h4 : 3'h0; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_265 = _decoded_signals_T_99 ? 3'h0 : _decoded_signals_T_264; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_266 = _decoded_signals_T_97 ? 3'h0 : _decoded_signals_T_265; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_267 = _decoded_signals_T_95 ? 3'h0 : _decoded_signals_T_266; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_268 = _decoded_signals_T_93 ? 3'h0 : _decoded_signals_T_267; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_269 = _decoded_signals_T_91 ? 3'h0 : _decoded_signals_T_268; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_270 = _decoded_signals_T_89 ? 3'h0 : _decoded_signals_T_269; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_271 = _decoded_signals_T_87 ? 3'h0 : _decoded_signals_T_270; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_272 = _decoded_signals_T_85 ? 3'h3 : _decoded_signals_T_271; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_273 = _decoded_signals_T_83 ? 3'h3 : _decoded_signals_T_272; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_274 = _decoded_signals_T_81 ? 3'h3 : _decoded_signals_T_273; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_275 = _decoded_signals_T_79 ? 3'h3 : _decoded_signals_T_274; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_276 = _decoded_signals_T_77 ? 3'h2 : _decoded_signals_T_275; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_277 = _decoded_signals_T_75 ? 3'h2 : _decoded_signals_T_276; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_278 = _decoded_signals_T_73 ? 3'h2 : _decoded_signals_T_277; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_279 = _decoded_signals_T_71 ? 3'h2 : _decoded_signals_T_278; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_280 = _decoded_signals_T_69 ? 3'h2 : _decoded_signals_T_279; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_281 = _decoded_signals_T_67 ? 3'h2 : _decoded_signals_T_280; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_282 = _decoded_signals_T_65 ? 3'h2 : _decoded_signals_T_281; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_283 = _decoded_signals_T_63 ? 3'h2 : _decoded_signals_T_282; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_284 = _decoded_signals_T_61 ? 3'h2 : _decoded_signals_T_283; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_285 = _decoded_signals_T_59 ? 3'h2 : _decoded_signals_T_284; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_286 = _decoded_signals_T_57 ? 3'h2 : _decoded_signals_T_285; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_287 = _decoded_signals_T_55 ? 3'h2 : _decoded_signals_T_286; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_288 = _decoded_signals_T_53 ? 3'h2 : _decoded_signals_T_287; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_289 = _decoded_signals_T_51 ? 3'h2 : _decoded_signals_T_288; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_290 = _decoded_signals_T_49 ? 3'h2 : _decoded_signals_T_289; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_291 = _decoded_signals_T_47 ? 3'h2 : _decoded_signals_T_290; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_292 = _decoded_signals_T_45 ? 3'h2 : _decoded_signals_T_291; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_293 = _decoded_signals_T_43 ? 3'h2 : _decoded_signals_T_292; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_294 = _decoded_signals_T_41 ? 3'h2 : _decoded_signals_T_293; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_295 = _decoded_signals_T_39 ? 3'h2 : _decoded_signals_T_294; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_296 = _decoded_signals_T_37 ? 3'h1 : _decoded_signals_T_295; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_297 = _decoded_signals_T_35 ? 3'h1 : _decoded_signals_T_296; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_298 = _decoded_signals_T_33 ? 3'h1 : _decoded_signals_T_297; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_299 = _decoded_signals_T_31 ? 3'h1 : _decoded_signals_T_298; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_300 = _decoded_signals_T_29 ? 3'h1 : _decoded_signals_T_299; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_301 = _decoded_signals_T_27 ? 3'h1 : _decoded_signals_T_300; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_302 = _decoded_signals_T_25 ? 3'h1 : _decoded_signals_T_301; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_303 = _decoded_signals_T_23 ? 3'h1 : _decoded_signals_T_302; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_304 = _decoded_signals_T_21 ? 3'h1 : _decoded_signals_T_303; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_305 = _decoded_signals_T_19 ? 3'h1 : _decoded_signals_T_304; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_306 = _decoded_signals_T_17 ? 3'h1 : _decoded_signals_T_305; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_307 = _decoded_signals_T_15 ? 3'h1 : _decoded_signals_T_306; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_308 = _decoded_signals_T_13 ? 3'h1 : _decoded_signals_T_307; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_309 = _decoded_signals_T_11 ? 3'h1 : _decoded_signals_T_308; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_310 = _decoded_signals_T_9 ? 3'h1 : _decoded_signals_T_309; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_311 = _decoded_signals_T_7 ? 3'h1 : _decoded_signals_T_310; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_312 = _decoded_signals_T_5 ? 3'h1 : _decoded_signals_T_311; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_313 = _decoded_signals_T_3 ? 3'h1 : _decoded_signals_T_312; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_316 = _decoded_signals_T_101 ? 4'h1 : 4'h0; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_317 = _decoded_signals_T_99 ? 4'h1 : _decoded_signals_T_316; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_318 = _decoded_signals_T_97 ? 4'h0 : _decoded_signals_T_317; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_319 = _decoded_signals_T_95 ? 4'h0 : _decoded_signals_T_318; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_320 = _decoded_signals_T_93 ? 4'h0 : _decoded_signals_T_319; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_321 = _decoded_signals_T_91 ? 4'h0 : _decoded_signals_T_320; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_322 = _decoded_signals_T_89 ? 4'h0 : _decoded_signals_T_321; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_323 = _decoded_signals_T_87 ? 4'h0 : _decoded_signals_T_322; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_324 = _decoded_signals_T_85 ? 4'h1 : _decoded_signals_T_323; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_325 = _decoded_signals_T_83 ? 4'h1 : _decoded_signals_T_324; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_326 = _decoded_signals_T_81 ? 4'h1 : _decoded_signals_T_325; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_327 = _decoded_signals_T_79 ? 4'h1 : _decoded_signals_T_326; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_328 = _decoded_signals_T_77 ? 4'hd : _decoded_signals_T_327; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_329 = _decoded_signals_T_75 ? 4'h0 : _decoded_signals_T_328; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_330 = _decoded_signals_T_73 ? 4'hb : _decoded_signals_T_329; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_331 = _decoded_signals_T_71 ? 4'ha : _decoded_signals_T_330; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_332 = _decoded_signals_T_69 ? 4'h9 : _decoded_signals_T_331; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_333 = _decoded_signals_T_67 ? 4'h8 : _decoded_signals_T_332; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_334 = _decoded_signals_T_65 ? 4'h8 : _decoded_signals_T_333; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_335 = _decoded_signals_T_63 ? 4'h7 : _decoded_signals_T_334; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_336 = _decoded_signals_T_61 ? 4'h7 : _decoded_signals_T_335; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_337 = _decoded_signals_T_59 ? 4'h6 : _decoded_signals_T_336; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_338 = _decoded_signals_T_57 ? 4'h6 : _decoded_signals_T_337; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_339 = _decoded_signals_T_55 ? 4'h1 : _decoded_signals_T_338; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_340 = _decoded_signals_T_53 ? 4'h1 : _decoded_signals_T_339; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_341 = _decoded_signals_T_51 ? 4'h1 : _decoded_signals_T_340; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_342 = _decoded_signals_T_49 ? 4'h1 : _decoded_signals_T_341; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_343 = _decoded_signals_T_47 ? 4'h1 : _decoded_signals_T_342; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_344 = _decoded_signals_T_45 ? 4'h1 : _decoded_signals_T_343; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_345 = _decoded_signals_T_43 ? 4'h1 : _decoded_signals_T_344; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_346 = _decoded_signals_T_41 ? 4'h1 : _decoded_signals_T_345; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_347 = _decoded_signals_T_39 ? 4'h1 : _decoded_signals_T_346; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_348 = _decoded_signals_T_37 ? 4'hd : _decoded_signals_T_347; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_349 = _decoded_signals_T_35 ? 4'hc : _decoded_signals_T_348; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_350 = _decoded_signals_T_33 ? 4'hb : _decoded_signals_T_349; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_351 = _decoded_signals_T_31 ? 4'ha : _decoded_signals_T_350; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_352 = _decoded_signals_T_29 ? 4'h9 : _decoded_signals_T_351; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_353 = _decoded_signals_T_27 ? 4'h8 : _decoded_signals_T_352; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_354 = _decoded_signals_T_25 ? 4'h7 : _decoded_signals_T_353; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_355 = _decoded_signals_T_23 ? 4'h6 : _decoded_signals_T_354; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_356 = _decoded_signals_T_21 ? 4'h6 : _decoded_signals_T_355; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_357 = _decoded_signals_T_19 ? 4'h5 : _decoded_signals_T_356; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_358 = _decoded_signals_T_17 ? 4'h4 : _decoded_signals_T_357; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_359 = _decoded_signals_T_15 ? 4'h4 : _decoded_signals_T_358; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_360 = _decoded_signals_T_13 ? 4'h4 : _decoded_signals_T_359; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_361 = _decoded_signals_T_11 ? 4'h3 : _decoded_signals_T_360; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_362 = _decoded_signals_T_9 ? 4'h3 : _decoded_signals_T_361; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_363 = _decoded_signals_T_7 ? 4'h2 : _decoded_signals_T_362; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_364 = _decoded_signals_T_5 ? 4'h2 : _decoded_signals_T_363; // @[Lookup.scala 34:39]
  wire [3:0] _decoded_signals_T_365 = _decoded_signals_T_3 ? 4'h1 : _decoded_signals_T_364; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_367 = _decoded_signals_T_103 ? 2'h2 : 2'h0; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_368 = _decoded_signals_T_101 ? 2'h0 : _decoded_signals_T_367; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_369 = _decoded_signals_T_99 ? 2'h0 : _decoded_signals_T_368; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_370 = _decoded_signals_T_97 ? 2'h0 : _decoded_signals_T_369; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_371 = _decoded_signals_T_95 ? 2'h0 : _decoded_signals_T_370; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_372 = _decoded_signals_T_93 ? 2'h0 : _decoded_signals_T_371; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_373 = _decoded_signals_T_91 ? 2'h0 : _decoded_signals_T_372; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_374 = _decoded_signals_T_89 ? 2'h0 : _decoded_signals_T_373; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_375 = _decoded_signals_T_87 ? 2'h0 : _decoded_signals_T_374; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_376 = _decoded_signals_T_85 ? 2'h0 : _decoded_signals_T_375; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_377 = _decoded_signals_T_83 ? 2'h0 : _decoded_signals_T_376; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_378 = _decoded_signals_T_81 ? 2'h0 : _decoded_signals_T_377; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_379 = _decoded_signals_T_79 ? 2'h0 : _decoded_signals_T_378; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_380 = _decoded_signals_T_77 ? 2'h0 : _decoded_signals_T_379; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_381 = _decoded_signals_T_75 ? 2'h2 : _decoded_signals_T_380; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_382 = _decoded_signals_T_73 ? 2'h0 : _decoded_signals_T_381; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_383 = _decoded_signals_T_71 ? 2'h0 : _decoded_signals_T_382; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_384 = _decoded_signals_T_69 ? 2'h0 : _decoded_signals_T_383; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_385 = _decoded_signals_T_67 ? 2'h0 : _decoded_signals_T_384; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_386 = _decoded_signals_T_65 ? 2'h0 : _decoded_signals_T_385; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_387 = _decoded_signals_T_63 ? 2'h0 : _decoded_signals_T_386; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_388 = _decoded_signals_T_61 ? 2'h0 : _decoded_signals_T_387; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_389 = _decoded_signals_T_59 ? 2'h0 : _decoded_signals_T_388; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_390 = _decoded_signals_T_57 ? 2'h0 : _decoded_signals_T_389; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_391 = _decoded_signals_T_55 ? 2'h0 : _decoded_signals_T_390; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_392 = _decoded_signals_T_53 ? 2'h0 : _decoded_signals_T_391; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_393 = _decoded_signals_T_51 ? 2'h1 : _decoded_signals_T_392; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_394 = _decoded_signals_T_49 ? 2'h1 : _decoded_signals_T_393; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_395 = _decoded_signals_T_47 ? 2'h1 : _decoded_signals_T_394; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_396 = _decoded_signals_T_45 ? 2'h1 : _decoded_signals_T_395; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_397 = _decoded_signals_T_43 ? 2'h1 : _decoded_signals_T_396; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_398 = _decoded_signals_T_41 ? 2'h1 : _decoded_signals_T_397; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_399 = _decoded_signals_T_39 ? 2'h1 : _decoded_signals_T_398; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_400 = _decoded_signals_T_37 ? 2'h0 : _decoded_signals_T_399; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_401 = _decoded_signals_T_35 ? 2'h0 : _decoded_signals_T_400; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_402 = _decoded_signals_T_33 ? 2'h0 : _decoded_signals_T_401; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_403 = _decoded_signals_T_31 ? 2'h0 : _decoded_signals_T_402; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_404 = _decoded_signals_T_29 ? 2'h0 : _decoded_signals_T_403; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_405 = _decoded_signals_T_27 ? 2'h0 : _decoded_signals_T_404; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_406 = _decoded_signals_T_25 ? 2'h0 : _decoded_signals_T_405; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_407 = _decoded_signals_T_23 ? 2'h0 : _decoded_signals_T_406; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_408 = _decoded_signals_T_21 ? 2'h0 : _decoded_signals_T_407; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_409 = _decoded_signals_T_19 ? 2'h0 : _decoded_signals_T_408; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_410 = _decoded_signals_T_17 ? 2'h0 : _decoded_signals_T_409; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_411 = _decoded_signals_T_15 ? 2'h0 : _decoded_signals_T_410; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_412 = _decoded_signals_T_13 ? 2'h0 : _decoded_signals_T_411; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_413 = _decoded_signals_T_11 ? 2'h0 : _decoded_signals_T_412; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_414 = _decoded_signals_T_9 ? 2'h0 : _decoded_signals_T_413; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_415 = _decoded_signals_T_7 ? 2'h0 : _decoded_signals_T_414; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_416 = _decoded_signals_T_5 ? 2'h0 : _decoded_signals_T_415; // @[Lookup.scala 34:39]
  wire [1:0] _decoded_signals_T_417 = _decoded_signals_T_3 ? 2'h0 : _decoded_signals_T_416; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_422 = _decoded_signals_T_97 ? 1'h0 : _decoded_signals_T_99 | (_decoded_signals_T_101 |
    _decoded_signals_T_103); // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_423 = _decoded_signals_T_95 ? 1'h0 : _decoded_signals_T_422; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_424 = _decoded_signals_T_93 ? 1'h0 : _decoded_signals_T_423; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_425 = _decoded_signals_T_91 ? 1'h0 : _decoded_signals_T_424; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_426 = _decoded_signals_T_89 ? 1'h0 : _decoded_signals_T_425; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_427 = _decoded_signals_T_87 ? 1'h0 : _decoded_signals_T_426; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_428 = _decoded_signals_T_85 ? 1'h0 : _decoded_signals_T_427; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_429 = _decoded_signals_T_83 ? 1'h0 : _decoded_signals_T_428; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_430 = _decoded_signals_T_81 ? 1'h0 : _decoded_signals_T_429; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_431 = _decoded_signals_T_79 ? 1'h0 : _decoded_signals_T_430; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_461 = _decoded_signals_T_19 | (_decoded_signals_T_21 | (_decoded_signals_T_23 | (
    _decoded_signals_T_25 | (_decoded_signals_T_27 | (_decoded_signals_T_29 | (_decoded_signals_T_31 | (
    _decoded_signals_T_33 | (_decoded_signals_T_35 | (_decoded_signals_T_37 | (_decoded_signals_T_39 | (
    _decoded_signals_T_41 | (_decoded_signals_T_43 | (_decoded_signals_T_45 | (_decoded_signals_T_47 | (
    _decoded_signals_T_49 | (_decoded_signals_T_51 | (_decoded_signals_T_53 | (_decoded_signals_T_55 | (
    _decoded_signals_T_57 | (_decoded_signals_T_59 | (_decoded_signals_T_61 | (_decoded_signals_T_63 | (
    _decoded_signals_T_65 | (_decoded_signals_T_67 | (_decoded_signals_T_69 | (_decoded_signals_T_71 | (
    _decoded_signals_T_73 | (_decoded_signals_T_75 | (_decoded_signals_T_77 | _decoded_signals_T_431))))))))))))))))))))
    ))))))))); // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_484 = _decoded_signals_T_77 ? 1'h0 : _decoded_signals_T_79 | (_decoded_signals_T_81 | (
    _decoded_signals_T_83 | _decoded_signals_T_85)); // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_485 = _decoded_signals_T_75 ? 1'h0 : _decoded_signals_T_484; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_486 = _decoded_signals_T_73 ? 1'h0 : _decoded_signals_T_485; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_487 = _decoded_signals_T_71 ? 1'h0 : _decoded_signals_T_486; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_488 = _decoded_signals_T_69 ? 1'h0 : _decoded_signals_T_487; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_489 = _decoded_signals_T_67 ? 1'h0 : _decoded_signals_T_488; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_490 = _decoded_signals_T_65 ? 1'h0 : _decoded_signals_T_489; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_491 = _decoded_signals_T_63 ? 1'h0 : _decoded_signals_T_490; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_492 = _decoded_signals_T_61 ? 1'h0 : _decoded_signals_T_491; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_493 = _decoded_signals_T_59 ? 1'h0 : _decoded_signals_T_492; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_494 = _decoded_signals_T_57 ? 1'h0 : _decoded_signals_T_493; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_495 = _decoded_signals_T_55 ? 1'h0 : _decoded_signals_T_494; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_496 = _decoded_signals_T_53 ? 1'h0 : _decoded_signals_T_495; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_497 = _decoded_signals_T_51 ? 1'h0 : _decoded_signals_T_496; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_498 = _decoded_signals_T_49 ? 1'h0 : _decoded_signals_T_497; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_499 = _decoded_signals_T_47 ? 1'h0 : _decoded_signals_T_498; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_500 = _decoded_signals_T_45 ? 1'h0 : _decoded_signals_T_499; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_501 = _decoded_signals_T_43 ? 1'h0 : _decoded_signals_T_500; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_502 = _decoded_signals_T_41 ? 1'h0 : _decoded_signals_T_501; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_503 = _decoded_signals_T_39 ? 1'h0 : _decoded_signals_T_502; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_504 = _decoded_signals_T_37 ? 1'h0 : _decoded_signals_T_503; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_505 = _decoded_signals_T_35 ? 1'h0 : _decoded_signals_T_504; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_506 = _decoded_signals_T_33 ? 1'h0 : _decoded_signals_T_505; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_507 = _decoded_signals_T_31 ? 1'h0 : _decoded_signals_T_506; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_508 = _decoded_signals_T_29 ? 1'h0 : _decoded_signals_T_507; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_509 = _decoded_signals_T_27 ? 1'h0 : _decoded_signals_T_508; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_510 = _decoded_signals_T_25 ? 1'h0 : _decoded_signals_T_509; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_511 = _decoded_signals_T_23 ? 1'h0 : _decoded_signals_T_510; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_512 = _decoded_signals_T_21 ? 1'h0 : _decoded_signals_T_511; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_513 = _decoded_signals_T_19 ? 1'h0 : _decoded_signals_T_512; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_514 = _decoded_signals_T_17 ? 1'h0 : _decoded_signals_T_513; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_515 = _decoded_signals_T_15 ? 1'h0 : _decoded_signals_T_514; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_516 = _decoded_signals_T_13 ? 1'h0 : _decoded_signals_T_515; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_517 = _decoded_signals_T_11 ? 1'h0 : _decoded_signals_T_516; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_518 = _decoded_signals_T_9 ? 1'h0 : _decoded_signals_T_517; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_519 = _decoded_signals_T_7 ? 1'h0 : _decoded_signals_T_518; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_520 = _decoded_signals_T_5 ? 1'h0 : _decoded_signals_T_519; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_521 = _decoded_signals_T_3 ? 1'h0 : _decoded_signals_T_520; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_532 = _decoded_signals_T_85 ? 3'h0 : 3'h6; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_533 = _decoded_signals_T_83 ? 3'h2 : _decoded_signals_T_532; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_534 = _decoded_signals_T_81 ? 3'h4 : _decoded_signals_T_533; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_535 = _decoded_signals_T_79 ? 3'h6 : _decoded_signals_T_534; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_536 = _decoded_signals_T_77 ? 3'h6 : _decoded_signals_T_535; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_537 = _decoded_signals_T_75 ? 3'h6 : _decoded_signals_T_536; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_538 = _decoded_signals_T_73 ? 3'h6 : _decoded_signals_T_537; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_539 = _decoded_signals_T_71 ? 3'h6 : _decoded_signals_T_538; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_540 = _decoded_signals_T_69 ? 3'h6 : _decoded_signals_T_539; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_541 = _decoded_signals_T_67 ? 3'h6 : _decoded_signals_T_540; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_542 = _decoded_signals_T_65 ? 3'h6 : _decoded_signals_T_541; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_543 = _decoded_signals_T_63 ? 3'h6 : _decoded_signals_T_542; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_544 = _decoded_signals_T_61 ? 3'h6 : _decoded_signals_T_543; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_545 = _decoded_signals_T_59 ? 3'h6 : _decoded_signals_T_544; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_546 = _decoded_signals_T_57 ? 3'h6 : _decoded_signals_T_545; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_547 = _decoded_signals_T_55 ? 3'h6 : _decoded_signals_T_546; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_548 = _decoded_signals_T_53 ? 3'h6 : _decoded_signals_T_547; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_549 = _decoded_signals_T_51 ? 3'h1 : _decoded_signals_T_548; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_550 = _decoded_signals_T_49 ? 3'h0 : _decoded_signals_T_549; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_551 = _decoded_signals_T_47 ? 3'h3 : _decoded_signals_T_550; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_552 = _decoded_signals_T_45 ? 3'h2 : _decoded_signals_T_551; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_553 = _decoded_signals_T_43 ? 3'h5 : _decoded_signals_T_552; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_554 = _decoded_signals_T_41 ? 3'h4 : _decoded_signals_T_553; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_555 = _decoded_signals_T_39 ? 3'h6 : _decoded_signals_T_554; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_556 = _decoded_signals_T_37 ? 3'h6 : _decoded_signals_T_555; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_557 = _decoded_signals_T_35 ? 3'h6 : _decoded_signals_T_556; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_558 = _decoded_signals_T_33 ? 3'h6 : _decoded_signals_T_557; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_559 = _decoded_signals_T_31 ? 3'h6 : _decoded_signals_T_558; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_560 = _decoded_signals_T_29 ? 3'h6 : _decoded_signals_T_559; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_561 = _decoded_signals_T_27 ? 3'h6 : _decoded_signals_T_560; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_562 = _decoded_signals_T_25 ? 3'h6 : _decoded_signals_T_561; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_563 = _decoded_signals_T_23 ? 3'h6 : _decoded_signals_T_562; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_564 = _decoded_signals_T_21 ? 3'h6 : _decoded_signals_T_563; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_565 = _decoded_signals_T_19 ? 3'h6 : _decoded_signals_T_564; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_566 = _decoded_signals_T_17 ? 3'h6 : _decoded_signals_T_565; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_567 = _decoded_signals_T_15 ? 3'h6 : _decoded_signals_T_566; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_568 = _decoded_signals_T_13 ? 3'h6 : _decoded_signals_T_567; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_569 = _decoded_signals_T_11 ? 3'h6 : _decoded_signals_T_568; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_570 = _decoded_signals_T_9 ? 3'h6 : _decoded_signals_T_569; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_571 = _decoded_signals_T_7 ? 3'h6 : _decoded_signals_T_570; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_572 = _decoded_signals_T_5 ? 3'h6 : _decoded_signals_T_571; // @[Lookup.scala 34:39]
  wire [2:0] _decoded_signals_T_573 = _decoded_signals_T_3 ? 3'h6 : _decoded_signals_T_572; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_578 = _decoded_signals_T_97 ? 1'h0 : _decoded_signals_T_99; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_579 = _decoded_signals_T_95 ? 1'h0 : _decoded_signals_T_578; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_580 = _decoded_signals_T_93 ? 1'h0 : _decoded_signals_T_579; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_581 = _decoded_signals_T_91 ? 1'h0 : _decoded_signals_T_580; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_582 = _decoded_signals_T_89 ? 1'h0 : _decoded_signals_T_581; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_583 = _decoded_signals_T_87 ? 1'h0 : _decoded_signals_T_582; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_584 = _decoded_signals_T_85 ? 1'h0 : _decoded_signals_T_583; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_585 = _decoded_signals_T_83 ? 1'h0 : _decoded_signals_T_584; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_586 = _decoded_signals_T_81 ? 1'h0 : _decoded_signals_T_585; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_587 = _decoded_signals_T_79 ? 1'h0 : _decoded_signals_T_586; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_588 = _decoded_signals_T_77 ? 1'h0 : _decoded_signals_T_587; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_589 = _decoded_signals_T_75 ? 1'h0 : _decoded_signals_T_588; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_590 = _decoded_signals_T_73 ? 1'h0 : _decoded_signals_T_589; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_591 = _decoded_signals_T_71 ? 1'h0 : _decoded_signals_T_590; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_592 = _decoded_signals_T_69 ? 1'h0 : _decoded_signals_T_591; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_594 = _decoded_signals_T_65 ? 1'h0 : _decoded_signals_T_67 | _decoded_signals_T_592; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_596 = _decoded_signals_T_61 ? 1'h0 : _decoded_signals_T_63 | _decoded_signals_T_594; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_598 = _decoded_signals_T_57 ? 1'h0 : _decoded_signals_T_59 | _decoded_signals_T_596; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_600 = _decoded_signals_T_53 ? 1'h0 : _decoded_signals_T_55 | _decoded_signals_T_598; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_601 = _decoded_signals_T_51 ? 1'h0 : _decoded_signals_T_600; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_602 = _decoded_signals_T_49 ? 1'h0 : _decoded_signals_T_601; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_603 = _decoded_signals_T_47 ? 1'h0 : _decoded_signals_T_602; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_604 = _decoded_signals_T_45 ? 1'h0 : _decoded_signals_T_603; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_605 = _decoded_signals_T_43 ? 1'h0 : _decoded_signals_T_604; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_606 = _decoded_signals_T_41 ? 1'h0 : _decoded_signals_T_605; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_607 = _decoded_signals_T_39 ? 1'h0 : _decoded_signals_T_606; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_608 = _decoded_signals_T_37 ? 1'h0 : _decoded_signals_T_607; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_609 = _decoded_signals_T_35 ? 1'h0 : _decoded_signals_T_608; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_610 = _decoded_signals_T_33 ? 1'h0 : _decoded_signals_T_609; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_611 = _decoded_signals_T_31 ? 1'h0 : _decoded_signals_T_610; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_612 = _decoded_signals_T_29 ? 1'h0 : _decoded_signals_T_611; // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_616 = _decoded_signals_T_21 ? 1'h0 : _decoded_signals_T_23 | (_decoded_signals_T_25 | (
    _decoded_signals_T_27 | _decoded_signals_T_612)); // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_619 = _decoded_signals_T_15 ? 1'h0 : _decoded_signals_T_17 | (_decoded_signals_T_19 |
    _decoded_signals_T_616); // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_622 = _decoded_signals_T_9 ? 1'h0 : _decoded_signals_T_11 | (_decoded_signals_T_13 |
    _decoded_signals_T_619); // @[Lookup.scala 34:39]
  wire  _decoded_signals_T_624 = _decoded_signals_T_5 ? 1'h0 : _decoded_signals_T_7 | _decoded_signals_T_622; // @[Lookup.scala 34:39]
  wire [2:0] _io_idu_to_exu_pc_sel_T = io_idu_to_exu_br_eq ? 3'h1 : 3'h0; // @[IDU.scala 115:20]
  wire [2:0] _io_idu_to_exu_pc_sel_T_2 = ~io_idu_to_exu_br_eq ? 3'h1 : 3'h0; // @[IDU.scala 116:20]
  wire [2:0] _io_idu_to_exu_pc_sel_T_4 = ~io_idu_to_exu_br_lt ? 3'h1 : 3'h0; // @[IDU.scala 117:20]
  wire [2:0] _io_idu_to_exu_pc_sel_T_6 = ~io_idu_to_exu_br_ltu ? 3'h1 : 3'h0; // @[IDU.scala 118:20]
  wire [2:0] _io_idu_to_exu_pc_sel_T_7 = io_idu_to_exu_br_lt ? 3'h1 : 3'h0; // @[IDU.scala 119:20]
  wire [2:0] _io_idu_to_exu_pc_sel_T_8 = io_idu_to_exu_br_ltu ? 3'h1 : 3'h0; // @[IDU.scala 120:20]
  wire [2:0] _io_idu_to_exu_pc_sel_T_10 = 4'h0 == br_type ? 3'h0 : 3'h4; // @[Mux.scala 81:58]
  wire [2:0] _io_idu_to_exu_pc_sel_T_12 = 4'h7 == br_type ? 3'h2 : _io_idu_to_exu_pc_sel_T_10; // @[Mux.scala 81:58]
  wire [2:0] _io_idu_to_exu_pc_sel_T_14 = 4'h8 == br_type ? 3'h3 : _io_idu_to_exu_pc_sel_T_12; // @[Mux.scala 81:58]
  wire [2:0] _io_idu_to_exu_pc_sel_T_16 = 4'h2 == br_type ? _io_idu_to_exu_pc_sel_T : _io_idu_to_exu_pc_sel_T_14; // @[Mux.scala 81:58]
  wire [2:0] _io_idu_to_exu_pc_sel_T_18 = 4'h1 == br_type ? _io_idu_to_exu_pc_sel_T_2 : _io_idu_to_exu_pc_sel_T_16; // @[Mux.scala 81:58]
  wire [2:0] _io_idu_to_exu_pc_sel_T_20 = 4'h3 == br_type ? _io_idu_to_exu_pc_sel_T_4 : _io_idu_to_exu_pc_sel_T_18; // @[Mux.scala 81:58]
  wire [2:0] _io_idu_to_exu_pc_sel_T_22 = 4'h4 == br_type ? _io_idu_to_exu_pc_sel_T_6 : _io_idu_to_exu_pc_sel_T_20; // @[Mux.scala 81:58]
  wire [2:0] _io_idu_to_exu_pc_sel_T_24 = 4'h5 == br_type ? _io_idu_to_exu_pc_sel_T_7 : _io_idu_to_exu_pc_sel_T_22; // @[Mux.scala 81:58]
  wire [2:0] _io_idu_to_exu_pc_sel_T_26 = 4'h6 == br_type ? _io_idu_to_exu_pc_sel_T_8 : _io_idu_to_exu_pc_sel_T_24; // @[Mux.scala 81:58]
  assign io_idu_to_exu_pc_sel = {{1'd0}, _io_idu_to_exu_pc_sel_T_26}; // @[IDU.scala 109:25]
  assign io_idu_to_exu_op1_sel = _decoded_signals_T_1 ? 2'h1 : _decoded_signals_T_261; // @[Lookup.scala 34:39]
  assign io_idu_to_exu_op2_sel = _decoded_signals_T_1 ? 3'h1 : _decoded_signals_T_313; // @[Lookup.scala 34:39]
  assign io_idu_to_exu_alu_op = _decoded_signals_T_1 ? 4'h1 : _decoded_signals_T_365; // @[Lookup.scala 34:39]
  assign io_idu_to_exu_wb_sel = _decoded_signals_T_1 ? 2'h0 : _decoded_signals_T_417; // @[Lookup.scala 34:39]
  assign io_idu_to_exu_reg_wen = _decoded_signals_T_1 | (_decoded_signals_T_3 | (_decoded_signals_T_5 | (
    _decoded_signals_T_7 | (_decoded_signals_T_9 | (_decoded_signals_T_11 | (_decoded_signals_T_13 | (
    _decoded_signals_T_15 | (_decoded_signals_T_17 | _decoded_signals_T_461)))))))); // @[Lookup.scala 34:39]
  assign io_idu_to_exu_mem_msk_type = _decoded_signals_T_1 ? 3'h6 : _decoded_signals_T_573; // @[Lookup.scala 34:39]
  assign io_idu_to_exu_alu_msk_type = _decoded_signals_T_1 ? 1'h0 : _decoded_signals_T_3 | _decoded_signals_T_624; // @[Lookup.scala 34:39]
  assign io_isEbreak = 32'h100073 == io_inst; // @[IDU.scala 129:27]
  assign io_inv_inst = ~decoded_signals_0; // @[IDU.scala 130:18]
  assign io_isWriteMem = _decoded_signals_T_1 ? 1'h0 : _decoded_signals_T_521; // @[Lookup.scala 34:39]
endmodule
