`include "ysyx_22050039_instpat.v"
`include "ysyx_22050039_all_inst.v"

module ysyx_22050039_IDU #(XLEN = 64, INST_LEN = 32, NR_REG = 32, REG_SEL = 5) (
	input clk,
	input rst,
	input [INST_LEN-1:0] inst,
	input [XLEN-1:0] exec_result,
	output reg [XLEN-1:0] src1,
	output reg [XLEN-1:0] src2,
	output [`ysyx_22050039_FUNC_LEN-1:0] func,
	output pc_wen 
);

	import "DPI-C" function void set_gpr_ptr(input logic [XLEN-1:0] a []);
	initial set_gpr_ptr(regs);  // rf为通用寄存器的二维数组变量

	// submodule1 - registers_heap: generate GPRS x0-x31
	wire [XLEN-1:0] regs [NR_REG-1:0];
	wire [NR_REG-1:0] reg_each_wen; 
	wire reg_total_wen;  // no drive yet TODO: not decied whether necessary yet

	ysyx_22050039_Reg #(XLEN, 0) reg_zero (clk, rst, exec_result, regs[0], reg_total_wen & reg_each_wen[0]); 
	genvar i; 
	generate
		for(i = 1; i < NR_REG; i = i+1) begin
//			ysyx_22050039_Reg #(XLEN, 0) gen_gprs (clk, rst, exec_result, regs[i], reg_total_wen & reg_each_wen[i]);
			ysyx_22050039_Reg #(XLEN, 0) gen_gprs (clk, rst, exec_result, regs[i], reg_total_wen & reg_each_wen[i]);
		end
	endgenerate

	// submodule2 - instruction decoder: decode inst
	wire [6:0] opcode;
	wire [2:0] funct3;
	wire [REG_SEL-1:0] rd;
	wire [REG_SEL-1:0] rs1;
	wire [REG_SEL-1:0] rs2;
	wire [6:0] funct7;
	wire [19:0] imm;
	wire R, I, S, B, U, J; // only 1 of these will be high
	reg [7+3+3*REG_SEL+7+20+6+3+1+1-1:0] bundle;

	assign {opcode, funct3, rd, rs1, rs2, funct7, imm, R, I, S, B, U, J, func,
		pc_wen, reg_total_wen} = bundle;

//  INSTPAT("??????? ????? ????? 000 ????? 11000 11", beq    , B, s->dnpc = src1 == src2 ? s->pc + dest : s->snpc);
//  INSTPAT("??????? ????? ????? 001 ????? 11000 11", bne	   , B, s->dnpc = src1 != src2 ? s->pc + dest : s->snpc); 
//  INSTPAT("??????? ????? ????? 110 ????? 11000 11", bltu   , B, s->dnpc = src1 < src2 ? s->pc + dest : s->snpc);
//  INSTPAT("??????? ????? ????? 101 ????? 11000 11", bge    , B, s->dnpc = (sword_t)src1 >= (sword_t)src2 ? s->pc + dest : s->snpc);
//  INSTPAT("??????? ????? ????? 111 ????? 11000 11", bgeu   , B, s->dnpc = src1 >= src2 ? s->pc + dest : s->snpc);
//  INSTPAT("??????? ????? ????? 100 ????? 11000 11", blt    , B, s->dnpc = (sword_t)src1 < (sword_t)src2 ? s->pc + dest : s->snpc);
//	// I
//  INSTPAT("??????? ????? ????? 100 ????? 00100 11", xori   , I, R(dest) = src1 ^ src2;);
//  INSTPAT("??????? ????? ????? 011 ????? 00100 11", sltiu  , I, R(dest) = src1 < src2;);
//  INSTPAT("000000? ????? ????? 001 ????? 00100 11", slli   , I, R(dest) = ((src1) << ((src2) & shift_mask)));
//  INSTPAT("000000? ????? ????? 101 ????? 00100 11", srli   , I, R(dest) = ((src1) >> ((src2) & shift_mask)));
//  INSTPAT("010000? ????? ????? 101 ????? 00100 11", srai   , I, R(dest) = ((sword_t)(src1) >> ((src2) & shift_mask)));
//  INSTPAT("??????? ????? ????? 111 ????? 00100 11", andi   , I, R(dest) = src1 & src2;);
//  INSTPAT("??????? ????? ????? 110 ????? 00100 11", ori    , I, R(dest) = src1 | src2;);
//  INSTPAT("??????? ????? ????? 000 ????? 00110 11", addiw  , I, R(dest) = sext32to64((src1) + (src2)));
//  INSTPAT("0000000 ????? ????? 001 ????? 00110 11", slliw  , I, R(dest) = sext32to64((uint32_t)(src1) << ((src2) & 0x1f)));
//  INSTPAT("0000000 ????? ????? 101 ????? 00110 11", srliw  , I, R(dest) = sext32to64((uint32_t)(src1) >> ((src2) & 0x1f)));
//  INSTPAT("0100000 ????? ????? 101 ????? 00110 11", sraiw  , I, R(dest) = sext32to64((int32_t)(src1) >> ((src2) & 0x1f)));
//  INSTPAT("??????? ????? ????? 010 ????? 00000 11", lw     , I, R(dest) = (sword_t)(int32_t)Mr(src1 + src2, 4));
//  INSTPAT("??????? ????? ????? 110 ????? 00000 11", lwu    , I, R(dest) = Mr(src1 + src2, 4));
//  INSTPAT("??????? ????? ????? 001 ????? 00000 11", lh     , I, R(dest) = (sword_t)(int16_t)Mr(src1 + src2, 2));
//  INSTPAT("??????? ????? ????? 101 ????? 00000 11", lhu    , I, R(dest) = Mr(src1 + src2, 2));
//  INSTPAT("??????? ????? ????? 000 ????? 00000 11", lb     , I, R(dest) = (sword_t)(int8_t)Mr(src1 + src2, 1));
//  INSTPAT("??????? ????? ????? 100 ????? 00000 11", lbu    , I, R(dest) = Mr(src1 + src2, 1));
//	// R
//  INSTPAT("0000000 ????? ????? 000 ????? 01110 11", addw   , R, R(dest) = sext32to64((src1) + (src2)));
//  INSTPAT("0100000 ????? ????? 000 ????? 01110 11", subw   , R, R(dest) = sext32to64((src1) - (src2)));
//  INSTPAT("0000001 ????? ????? 000 ????? 01110 11", mulw   , R, R(dest) = sext32to64((src1) * (src2)));
//  INSTPAT("0000001 ????? ????? 100 ????? 01110 11", divw   , R, R(dest) = sext32to64((int32_t)(src1) / ( int32_t)(src2)));
//  INSTPAT("0000001 ????? ????? 101 ????? 01110 11", divuw  , R, R(dest) = sext32to64((uint32_t)(src1) / (uint32_t)(src2)));
//  INSTPAT("0000000 ????? ????? 001 ????? 01110 11", sllw   , R, R(dest) = sext32to64((uint32_t)(src1) << ((src2) & 0x1f)));
//  INSTPAT("0000000 ????? ????? 101 ????? 01110 11", srlw   , R, R(dest) = sext32to64((uint32_t)(src1) >> ((src2) & 0x1f)));
//  INSTPAT("0100000 ????? ????? 101 ????? 01110 11", sraw   , R, R(dest) = sext32to64((int32_t)(src1) >> ((src2) & 0x1f)));
//  INSTPAT("0000001 ????? ????? 110 ????? 01110 11", remw   , R, R(dest) = sext32to64((int32_t)(src1) % ( int32_t)(src2)));
//  INSTPAT("0000001 ????? ????? 111 ????? 01110 11", remuw  , R, R(dest) = sext32to64((uint32_t)(src1) % (uint32_t)(src2)));
//  INSTPAT("0100000 ????? ????? 000 ????? 01100 11", sub    , R, R(dest) = src1 - src2;);
//  INSTPAT("0000000 ????? ????? 110 ????? 01100 11", or     , R, R(dest) = src1 | src2;);
//  INSTPAT("0000000 ????? ????? 000 ????? 01100 11", add    , R, R(dest) = src1 + src2;);
//  INSTPAT("0000001 ????? ????? 000 ????? 01100 11", mul    , R, R(dest) = src1 * src2;);
//  INSTPAT("0000000 ????? ????? 100 ????? 01100 11", xor    , R, R(dest) = src1 ^ src2;);
//  INSTPAT("0000000 ????? ????? 001 ????? 01100 11", sll    , R, R(dest) = src1 << (src2 & shift_mask));
//  INSTPAT("0000000 ????? ????? 010 ????? 01100 11", slt    , R, R(dest) = (sword_t)src1 < (sword_t)src2;);
//  INSTPAT("0000000 ????? ????? 011 ????? 01100 11", sltu   , R, R(dest) = src1 < src2;);
//  INSTPAT("0000000 ????? ????? 111 ????? 01100 11", and    , R, R(dest) = src1 & src2;);
//  INSTPAT("0000001 ????? ????? 100 ????? 01100 11", div    , R, R(dest) = (sword_t)src1 / (sword_t)src2;);
//  INSTPAT("0000001 ????? ????? 101 ????? 01100 11", divu   , R, R(dest) = src1 / src2;);
//  INSTPAT("0000001 ????? ????? 110 ????? 01100 11", rem    , R, R(dest) = (sword_t)(src1) % (sword_t)(src2));
//  INSTPAT("0000001 ????? ????? 111 ????? 01100 11", remu   , R, R(dest) = src1 % src2;);
//	// S
//  INSTPAT("??????? ????? ????? 010 ????? 01000 11", sw     , S, Mw(src1 + dest, 4, src2));
//  INSTPAT("??????? ????? ????? 001 ????? 01000 11", sh     , S, Mw(src1 + dest, 2, src2));
//  INSTPAT("??????? ????? ????? 000 ????? 01000 11", sb     , S, Mw(src1 + dest, 1, src2));
//	// jmp
//
//  INSTPAT("??????? ????? ????? 011 ????? 00000 11", ld     , I, R(dest) = Mr(src1 + src2, 8));


	`ysyx_22050039_INSTPAT_START()
			// I-type
			`ysyx_22050039_INSTPAT(32'b?????????????????000?????0010011, {{8{inst[31]}}, inst[31:20]}, Itype, Addi, `ysyx_22050039_NO_WPC, `ysyx_22050039_WREG)
			`ysyx_22050039_INSTPAT(32'b?????????????????000?????1100111, {{8{inst[31]}}, inst[31:20]}, Itype, Jalr, `ysyx_22050039_WPC, `ysyx_22050039_WREG)
			// U-type
			`ysyx_22050039_INSTPAT(32'b?????????????????????????0010111, inst[31:12], Utype, Auipc, `ysyx_22050039_NO_WPC, `ysyx_22050039_WREG)
			`ysyx_22050039_INSTPAT(32'b?????????????????????????0110111, inst[31:12], Utype, Lui, `ysyx_22050039_NO_WPC, `ysyx_22050039_WREG)
			// S-type
			`ysyx_22050039_INSTPAT(32'b?????????????????011?????0100011, {{8{inst[31]}}, inst[31:25], inst[11:7]}, Stype, Sd, `ysyx_22050039_NO_WPC, `ysyx_22050039_NO_WREG)
			// J-type
			`ysyx_22050039_INSTPAT(32'b?????????????????????????1101111, {inst[31], inst[19:12], inst[20], inst[30:21]}, Jtype, Jal, `ysyx_22050039_WPC, `ysyx_22050039_WREG)
			// ebreak
			`ysyx_22050039_INSTPAT(32'b00000000000100000000000001110011, 20'b0, Special, Ebreak, `ysyx_22050039_NO_WPC, `ysyx_22050039_NO_WREG)
			// invalid
			`ysyx_22050039_INSTINVALID()
	`ysyx_22050039_INSTPAT_END()

	// submodule3 - define src1 src2 TODO: maybe we need to determine rd here
	// the future
	wire [5:0] inst_type;
	assign inst_type = {R, I, S, B, U, J};

	always@(*) begin	
		src1 = 0;
		src2 = 0;
		case(inst_type)
			// R
			Rtype		: begin src1 = regs[rs1]; src2 = regs[rs2]; end
			// I
			Itype		: begin src1 = regs[rs1]; src2 = {{44{imm[19]}}, imm}; end
			// S
			Stype		: ; // empty now
			// B
			Btype		: assert(0); // empty now
			// U
			Utype		: begin src1 = {{32{imm[19]}}, imm, 12'b0}; end
			// J
			Jtype		: begin src1 = {{43{imm[19]}}, imm, 1'b0}; end
			// ebreak and invalid
			Special	: ;	
			default : assert(0); 
		endcase
	end

	// submodule4 - reg addressing: 5-32 decoder 
	// Only 1 bit of output can be high, and that is the reg to write
	ysyx_22050039_MuxKey #(NR_REG, REG_SEL, NR_REG) selDestR (
		.out(reg_each_wen),
		.key(rd),
		.lut({
			5'd0, 32'h0000_0000, // $zero is always 0
			5'd1, 32'h0000_0002, 
			5'd2, 32'h0000_0004, 
			5'd3, 32'h0000_0008, 
			5'd4, 32'h0000_0010, 
			5'd5, 32'h0000_0020, 
			5'd6, 32'h0000_0040, 
			5'd7, 32'h0000_0080, 
			5'd8, 32'h0000_0100, 
			5'd9, 32'h0000_0200, 
			5'd10, 32'h0000_0400, 
			5'd11, 32'h0000_0800, 
			5'd12, 32'h0000_1000, 
			5'd13, 32'h0000_2000, 
			5'd14, 32'h0000_4000, 
			5'd15, 32'h0000_8000, 
			5'd16, 32'h0001_0000, 
			5'd17, 32'h0002_0000, 
			5'd18, 32'h0004_0000, 
			5'd19, 32'h0008_0000, 
			5'd20, 32'h0010_0000, 
			5'd21, 32'h0020_0000, 
			5'd22, 32'h0040_0000, 
			5'd23, 32'h0080_0000, 
			5'd24, 32'h0100_0000, 
			5'd25, 32'h0200_0000, 
			5'd26, 32'h0400_0000, 
			5'd27, 32'h0800_0000, 
			5'd28, 32'h1000_0000, 
			5'd29, 32'h2000_0000, 
			5'd30, 32'h4000_0000, 
			5'd31, 32'h8000_0000 
		})
	);

	always@(posedge clk) begin
		$display("inst_type = %d, func = %d, src1 = %x, src2 = %x", inst_type,
			func, src1, src2);
	end

endmodule

