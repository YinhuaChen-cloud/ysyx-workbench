`define INSTPAT_START() \
	always@(*) begin
	
`define INSTPAT_END() \
	end
