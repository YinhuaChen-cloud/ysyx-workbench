`define INSTPAT_START() \
	always@(*) begin
	
`define INSTPAT_END() \
	end

module ysyx_22050039_macro();
endmodule
