module ysyx_22050039_EXU
endmodule
