module ysyx_22050039_IDU
endmodule
