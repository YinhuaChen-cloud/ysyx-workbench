module ysyx_22050039_IFU(
	
);
	reg []

endmodule
